module risc ();

endmodule